library verilog;
use verilog.vl_types.all;
entity digital_circuits_final_work_vlg_vec_tst is
end digital_circuits_final_work_vlg_vec_tst;
